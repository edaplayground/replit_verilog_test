module test;

  initial
    $display("hello world!");

endmodule
